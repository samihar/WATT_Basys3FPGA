`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:07:48 06/12/2014 
// Design Name: 
// Module Name:    adder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder(
input [7:0] a,
input [7:0] b,
input clk,
input cin,
output reg [7:0] sum,
output reg [7:0] diff,
output reg cout

);
/*
YOUR CODE HERE
*/
endmodule

